

module square_demo (
    input clk,
    input [10:0] x, y,                // Current pixel coordinates (x and y)
    output [11:0] vga_rgb
);

// Internal signals


initial begin
    
end
reg [11:0] use_rgb;
initial  use_rgb = 0;
reg [3:0] r, g, b;                    // Individual RGB color channels

reg start;
reg [30:154] rowBuffer [30:110];
reg [155:346] numBuffer [30:110];
reg [15:0] numIt;
reg [15:0] statIt;
reg [15:0] thingIt;
reg [23:0] stats [7:0];
reg [10:0] currStat;
reg [40:0] count;
reg valid;
initial begin
    numIt = 30;
    statIt = 0;
    stats[0] = 24'h8;
    stats[1] = 24'h9;
    stats[2] = 24'ha;
    stats[3] = 24'hb;
    stats[4] = 24'hc;
    stats[5] = 24'hd;
    stats[6] = 24'he;
    stats[7] = 24'hf;
    currStat = 0;
    thingIt = 0;
    valid = 0;
    count = 0;
    
    rowBuffer[30] = 125'b00111000001110000111001111100011110001111001111100011110000000001111100011100011111000111000100000000000000000000000000;
    rowBuffer[31] = 125'b01000100010000001000001000000100000010000001000000100000000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[32] = 125'b01000100100000010000001000000100000010000001000000100000000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[33] = 125'b01111100100000010000001111100011100001110001111100011100000000000010000100010000100001111100100000000000000000000000000;
    rowBuffer[34] = 125'b01000100100000010000001000000000010000001001000000000010000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[35] = 125'b01000100010000001000001000000000010000001001000000000010000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[36] = 125'b01000100001110000111001111100111100011110001111100111100000000000010000011100000100001000100111110000000000000000000000;
    rowBuffer[37] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[38] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[39] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
    rowBuffer[40] = 125'b01000100111100011111001111100111110000000001000100111110011111000000000111110001110001111100011100010000000000000000000;
    rowBuffer[41] = 125'b01000100100010000100000010000100000000000001000100001000000100000000000001000010001000010000100010010000000111000000000;
    rowBuffer[42] = 125'b01000100100010000100000010000100000000000001000100001000000100000000000001000010001000010000100010010000000111000000000;
    rowBuffer[43] = 125'b01010100111100000100000010000111110000000001111100001000000100000000000001000010001000010000111110010000000000000000000;
    rowBuffer[44] = 125'b01010100101000000100000010000100000000000001000100001000000100000000000001000010001000010000100010010000000111000000000;
    rowBuffer[45] = 125'b01101100100100000100000010000100000000000001000100001000000100000000000001000010001000010000100010010000000111000000000;
    rowBuffer[46] = 125'b01000100100010011111000010000111110000000001000100111110000100000000000001000001110000010000100010011111000000000000000;
    rowBuffer[47] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[48] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[49] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
    rowBuffer[50] = 125'b01111000111110001110001111000000000010001001111100111110000000001111100011100011111000111000100000000000000000000000000;
    rowBuffer[51] = 125'b01000100100000010001001000100000000010001000010000001000000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[52] = 125'b01000100100000010001001000100000000010001000010000001000000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[53] = 125'b01111000111110011111001000100000000011111000010000001000000000000010000100010000100001111100100000000000000000000000000;
    rowBuffer[54] = 125'b01010000100000010001001000100000000010001000010000001000000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[55] = 125'b01001000100000010001001000100000000010001000010000001000000000000010000100010000100001000100100000001110000000000000000;
    rowBuffer[56] = 125'b01000100111110010001001111000000000010001001111100001000000000000010000011100000100001000100111110000000000000000000000;
    rowBuffer[57] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[58] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[59] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
    rowBuffer[60] = 125'b01000100111100011111001111100111110000000001000100111110001111000111100000000011111000111000111110001110001000000000000;
    rowBuffer[61] = 125'b01000100100010000100000010000100000000000001101100001000010000001000000000000000100001000100001000010001001000000011100;
    rowBuffer[62] = 125'b01000100100010000100000010000100000000000001010100001000010000001000000000000000100001000100001000010001001000000011100;
    rowBuffer[63] = 125'b01010100111100000100000010000111110000000001010100001000001110000111000000000000100001000100001000011111001000000000000;
    rowBuffer[64] = 125'b01010100101000000100000010000100000000000001000100001000000001000000100000000000100001000100001000010001001000000011100;
    rowBuffer[65] = 125'b01101100100100000100000010000100000000000001000100001000000001000000100000000000100001000100001000010001001000000011100;
    rowBuffer[66] = 125'b01000100100010011111000010000111110000000001000100111110011110001111000000000000100000111000001000010001001111100000000;
    rowBuffer[67] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[68] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[69] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
    rowBuffer[70] = 125'b01111000111110001110001111000000000010001001111100011110001111000000000111110001110001111100011100010000000000000000000;
    rowBuffer[71] = 125'b01000100100000010001001000100000000011011000010000100000010000000000000001000010001000010000100010010000000111000000000;
    rowBuffer[72] = 125'b01000100100000010001001000100000000010101000010000100000010000000000000001000010001000010000100010010000000111000000000;
    rowBuffer[73] = 125'b01111000111110011111001000100000000010101000010000011100001110000000000001000010001000010000111110010000000000000000000;
    rowBuffer[74] = 125'b01010000100000010001001000100000000010001000010000000010000001000000000001000010001000010000100010010000000111000000000;
    rowBuffer[75] = 125'b01001000100000010001001000100000000010001000010000000010000001000000000001000010001000010000100010010000000111000000000;
    rowBuffer[76] = 125'b01000100111110010001001111000000000010001001111100111100011110000000000001000001110000010000100010011111000000000000000;
    rowBuffer[77] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[78] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[79] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
    rowBuffer[80] = 125'b01111100100010001111001111100000000011111000111000111110001110001000000000000000000000000000000000000000000000000000000;
    rowBuffer[81] = 125'b00010000110010010000000010000000000000100001000100001000010001001000000011100000000000000000000000000000000000000000000;
    rowBuffer[82] = 125'b00010000101010010000000010000000000000100001000100001000010001001000000011100000000000000000000000000000000000000000000;
    rowBuffer[83] = 125'b00010000101010001110000010000000000000100001000100001000011111001000000000000000000000000000000000000000000000000000000;
    rowBuffer[84] = 125'b00010000100110000001000010000000000000100001000100001000010001001000000011100000000000000000000000000000000000000000000;
    rowBuffer[85] = 125'b00010000100010000001000010000000000000100001000100001000010001001000000011100000000000000000000000000000000000000000000;
    rowBuffer[86] = 125'b01111100100010011110000010000000000000100000111000001000010001001111100000000000000000000000000000000000000000000000000;
    rowBuffer[87] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[88] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[89] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
    rowBuffer[90] = 125'b01000100111110011111000000000111110001110001111100011100010000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[91] = 125'b01000100001000000100000000000001000010001000010000100010010000000111000000000000000000000000000000000000000000000000000;
    rowBuffer[92] = 125'b01000100001000000100000000000001000010001000010000100010010000000111000000000000000000000000000000000000000000000000000;
    rowBuffer[93] = 125'b01111100001000000100000000000001000010001000010000111110010000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[94] = 125'b01000100001000000100000000000001000010001000010000100010010000000111000000000000000000000000000000000000000000000000000;
    rowBuffer[95] = 125'b01000100001000000100000000000001000010001000010000100010010000000111000000000000000000000000000000000000000000000000000;
    rowBuffer[96] = 125'b01000100111110000100000000000001000001110000010000100010011111000000000000000000000000000000000000000000000000000000000;
    rowBuffer[97] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[98] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[99] = 125'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    
    rowBuffer[100] = 125'b0100010011111000111100011110000000001111100011100011111000111000100000000000000000000000000000000000000000000000000000;
    rowBuffer[101] = 125'b0110110000100001000000100000000000000010000100010000100001000100100000001110000000000000000000000000000000000000000000;
    rowBuffer[102] = 125'b0101010000100001000000100000000000000010000100010000100001000100100000001110000000000000000000000000000000000000000000;
    rowBuffer[103] = 125'b0101010000100000111000011100000000000010000100010000100001111100100000000000000000000000000000000000000000000000000000;
    rowBuffer[104] = 125'b0100010000100000000100000010000000000010000100010000100001000100100000001110000000000000000000000000000000000000000000;
    rowBuffer[105] = 125'b0100010000100000000100000010000000000010000100010000100001000100100000001110000000000000000000000000000000000000000000;
    rowBuffer[106] = 125'b0100010011111001111000111100000000000010000011100000100001000100111110000000000000000000000000000000000000000000000000;
    rowBuffer[107] = 125'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[108] = 125'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    rowBuffer[109] = 125'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;

    numBuffer[30] = 192'b0;
    numBuffer[31] = 192'b0;
    numBuffer[32] = 192'b0;
    numBuffer[33] = 192'b0;
    numBuffer[34] = 192'b0;
    numBuffer[35] = 192'b0;
    numBuffer[36] = 192'b0;
    numBuffer[37] = 192'b0;
    numBuffer[38] = 192'b0;
    numBuffer[39] = 192'b0;
    numBuffer[40] = 192'b0;
    numBuffer[41] = 192'b0;
    numBuffer[42] = 192'b0;
    numBuffer[43] = 192'b0;
    numBuffer[44] = 192'b0;
    numBuffer[45] = 192'b0;
    numBuffer[46] = 192'b0;
    numBuffer[47] = 192'b0;
    numBuffer[48] = 192'b0;
    numBuffer[49] = 192'b0;
    numBuffer[50] = 192'b0;
    numBuffer[51] = 192'b0;
    numBuffer[52] = 192'b0;
    numBuffer[53] = 192'b0;
    numBuffer[54] = 192'b0;
    numBuffer[55] = 192'b0;
    numBuffer[56] = 192'b0;
    numBuffer[57] = 192'b0;
    numBuffer[58] = 192'b0;
    numBuffer[59] = 192'b0;
    numBuffer[60] = 192'b0;
    numBuffer[61] = 192'b0;
    numBuffer[62] = 192'b0;
    numBuffer[63] = 192'b0;
    numBuffer[64] = 192'b0;
    numBuffer[65] = 192'b0;
    numBuffer[66] = 192'b0;
    numBuffer[67] = 192'b0;
    numBuffer[68] = 192'b0;
    numBuffer[69] = 192'b0;
    numBuffer[70] = 192'b0;
    numBuffer[71] = 192'b0;
    numBuffer[72] = 192'b0;
    numBuffer[73] = 192'b0;
    numBuffer[74] = 192'b0;
    numBuffer[75] = 192'b0;
    numBuffer[76] = 192'b0;
    numBuffer[77] = 192'b0;
    numBuffer[78] = 192'b0;
    numBuffer[79] = 192'b0;
    numBuffer[80] = 192'b0;
    numBuffer[81] = 192'b0;
    numBuffer[82] = 192'b0;
    numBuffer[83] = 192'b0;
    numBuffer[84] = 192'b0;
    numBuffer[85] = 192'b0;
    numBuffer[86] = 192'b0;
    numBuffer[87] = 192'b0;
    numBuffer[88] = 192'b0;
    numBuffer[89] = 192'b0;
    numBuffer[90] = 192'b0;
    numBuffer[91] = 192'b0;
    numBuffer[92] = 192'b0;
    numBuffer[93] = 192'b0;
    numBuffer[94] = 192'b0;
    numBuffer[95] = 192'b0;
    numBuffer[96] = 192'b0;
    numBuffer[97] = 192'b0;
    numBuffer[98] = 192'b0;
    numBuffer[99] = 192'b0;
    numBuffer[100] = 192'b0;
    numBuffer[101] = 192'b0;
    numBuffer[102] = 192'b0;
    numBuffer[103] = 192'b0;
    numBuffer[104] = 192'b0;
    numBuffer[105] = 192'b0;
    numBuffer[106] = 192'b0;
    numBuffer[107] = 192'b0;
    numBuffer[108] = 192'b0;
    numBuffer[109] = 192'b0;
end




// Combinational logic to set color based on pixel position
always @(posedge clk) begin
        r = use_rgb[3:0];
        g = use_rgb[7:4];
        b = use_rgb[11:8];
        if(y > 29 && y < 110) begin
            if(x > 29 && x < 155)begin
               if(rowBuffer[y][x])begin
                    r = 4'b1111 - use_rgb[3:0];
                    g = 4'b1111 - use_rgb[7:4];
                    b = 4'b1111 - use_rgb[11:8];
               end
            end
            else if(x > 154 && x < 347)begin
                if(numBuffer[y][x])begin
                    r = 4'b1111 - use_rgb[3:0];
                    g = 4'b1111 - use_rgb[7:4];
                    b = 4'b1111 - use_rgb[11:8];
               end
            end
        end
end

always @(posedge clk)begin
    count = count + 1;
    if(numIt < 110)begin
        if(statIt < 8)begin
                    case (stats[statIt][3:0])
                        4'b0000: begin
                            numBuffer[numIt][340:346] = 7'b0011100;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100010;
                            numBuffer[numIt+3][340:346] = 7'b0100010;
                            numBuffer[numIt+4][340:346] = 7'b0100010;
                            numBuffer[numIt+5][340:346] = 7'b0100010;
                            numBuffer[numIt+6][340:346] = 7'b0011100;
                        end
                        4'b0001: begin
                            numBuffer[numIt][340:346] = 7'b0011100;
                            numBuffer[numIt+1][340:346] = 7'b0011100;
                            numBuffer[numIt+2][340:346] = 7'b0011100;
                            numBuffer[numIt+3][340:346] = 7'b0011100;
                            numBuffer[numIt+4][340:346] = 7'b0011100;
                            numBuffer[numIt+5][340:346] = 7'b0011100;
                            numBuffer[numIt+6][340:346] = 7'b0011100;
                        end
                        4'b0010: begin
                            numBuffer[numIt][340:346] = 7'b0011100;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100110;
                            numBuffer[numIt+3][340:346] = 7'b0001100;
                            numBuffer[numIt+4][340:346] = 7'b0011000;
                            numBuffer[numIt+5][340:346] = 7'b0110000;
                            numBuffer[numIt+6][340:346] = 7'b0111110;
                        end
                        4'b0011: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt + 1][340:346] = 7'b0000010;
                            numBuffer[numIt + 2][340:346] = 7'b0000010;
                            numBuffer[numIt + 3][340:346] = 7'b0111110;
                            numBuffer[numIt + 4][340:346] = 7'b0000010;
                            numBuffer[numIt + 5][340:346] = 7'b0000010;
                            numBuffer[numIt + 6][340:346] = 7'b0111110;
                        end
                        4'b0100: begin
                            numBuffer[numIt][340:346] = 7'b0100010;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100010;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0000010;
                            numBuffer[numIt+5][340:346] = 7'b0000010;
                            numBuffer[numIt+6][340:346] = 7'b0000010;
                        end
                        4'b0101: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt+1][340:346] = 7'b0100000;
                            numBuffer[numIt+2][340:346] = 7'b0100000;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0000010;
                            numBuffer[numIt+5][340:346] = 7'b0000010;
                            numBuffer[numIt+6][340:346] = 7'b0111110;
                        end
                        4'b0110: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt+1][340:346] = 7'b0100000;
                            numBuffer[numIt+2][340:346] = 7'b0100000;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0100010;
                            numBuffer[numIt+5][340:346] = 7'b0100010;
                            numBuffer[numIt+6][340:346] = 7'b0111110;
                        end
                        4'b0111: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt+1][340:346] = 7'b0000010;
                            numBuffer[numIt+2][340:346] = 7'b0000100;
                            numBuffer[numIt+3][340:346] = 7'b0001000;
                            numBuffer[numIt+4][340:346] = 7'b0010000;
                            numBuffer[numIt+5][340:346] = 7'b0100000;
                            numBuffer[numIt+6][340:346] = 7'b0100000;
                        end
                        4'b1000: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100010;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0100010;
                            numBuffer[numIt+5][340:346] = 7'b0100010;
                            numBuffer[numIt+6][340:346] = 7'b0111110;
                        end
                        4'b1001: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100010;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0000010;
                            numBuffer[numIt+5][340:346] = 7'b0000010;
                            numBuffer[numIt+6][340:346] = 7'b0111110;
                        end
                        4'b1010: begin
                            numBuffer[numIt][340:346] = 7'b0011100;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100010;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0100010;
                            numBuffer[numIt+5][340:346] = 7'b0100010;
                            numBuffer[numIt+6][340:346] = 7'b0100010;
                        end
                        4'b1011: begin
                            numBuffer[numIt][340:346] = 7'b0111100;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100010;
                            numBuffer[numIt+3][340:346] = 7'b0111100;
                            numBuffer[numIt+4][340:346] = 7'b0100010;
                            numBuffer[numIt+5][340:346] = 7'b0100010;
                            numBuffer[numIt+6][340:346] = 7'b0111100;
                        end
                        4'b1100: begin
                            numBuffer[numIt][340:346] = 7'b0001110;
                            numBuffer[numIt+1][340:346] = 7'b0010000;
                            numBuffer[numIt+2][340:346] = 7'b0100000;
                            numBuffer[numIt+3][340:346] = 7'b0100000;
                            numBuffer[numIt+4][340:346] = 7'b0100000;
                            numBuffer[numIt+5][340:346] = 7'b0010000;
                            numBuffer[numIt+6][340:346] = 7'b0001110;
                        end
                        4'b1101: begin
                            numBuffer[numIt][340:346] = 7'b0111100;
                            numBuffer[numIt+1][340:346] = 7'b0100010;
                            numBuffer[numIt+2][340:346] = 7'b0100010;
                            numBuffer[numIt+3][340:346] = 7'b0100010;
                            numBuffer[numIt+4][340:346] = 7'b0100010;
                            numBuffer[numIt+5][340:346] = 7'b0100010;
                            numBuffer[numIt+6][340:346] = 7'b0111100;
                        end
                        4'b1110: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt+1][340:346] = 7'b0100000;
                            numBuffer[numIt+2][340:346] = 7'b0100000;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0100000;
                            numBuffer[numIt+5][340:346] = 7'b0100000;
                            numBuffer[numIt+6][340:346] = 7'b0111110;
                        end
                        4'b1111: begin
                            numBuffer[numIt][340:346] = 7'b0111110;
                            numBuffer[numIt+1][340:346] = 7'b0100000;
                            numBuffer[numIt+2][340:346] = 7'b0100000;
                            numBuffer[numIt+3][340:346] = 7'b0111110;
                            numBuffer[numIt+4][340:346] = 7'b0100000;
                            numBuffer[numIt+5][340:346] = 7'b0100000;
                            numBuffer[numIt+6][340:346] = 7'b0100000;
                        end
                        default: begin
                            numBuffer[numIt][340:346] = 7'b0000000;
                            numBuffer[numIt+1][340:346] = 7'b0000000;
                            numBuffer[numIt+2][340:346] = 7'b0000000;
                            numBuffer[numIt+3][340:346] = 7'b0000000;
                            numBuffer[numIt+4][340:346] = 7'b0000000;
                            numBuffer[numIt+5][340:346] = 7'b0000000;
                            numBuffer[numIt+6][340:346] = 7'b0000000;
                        end
                    endcase

                    statIt = statIt + 1;
                    numIt = numIt + 10;
            end
        //statIt = 0;
        
    end
    //numIt = 0;
end

// Output the final RGB value (reordered from {r,g,b} to {b,g,r})
assign vga_rgb = {b, g, r};   // Note: VGA often uses BGR order instead of RGB

endmodule